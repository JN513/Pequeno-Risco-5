module top (
    input clk25
);

always @(posedge clk25 ) begin

end

endmodule
