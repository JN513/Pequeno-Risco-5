module Control_Unit (
    input wire [6:0]instrution_opcode,
    output reg branch,
    output reg memory_read,
    output reg memory_to_reg,
    output reg [1:0] aluop,
    output reg memory_write,
    output reg alu_src,
    output reg reg_write
);

always @(*) begin
    case (instrution_opcode)
        7'b0110011: begin // R type instruction 
            alu_src = 0;
            memory_to_reg = 0;
            reg_write = 1;
            memory_read = 0;
            memory_write = 1;
            branch = 0;
            aluop = 2'b10;
        end

        7'b0000011: begin // lw instruction 
            alu_src = 1;
            memory_to_reg = 1;
            reg_write = 1;
            memory_read = 1;
            memory_write = 0;
            branch = 0;
            aluop = 2'b00;
        end

        7'b0100011: begin // sw instruction 
            alu_src = 1;
            memory_to_reg = x;
            reg_write = 0;
            memory_read = 0;
            memory_write = 1;
            branch = 0;
            aluop = 2'b00;
        end

        7'b1100011: begin // beq instruction 
            alu_src = 0;
            memory_to_reg = x;
            reg_write = 0;
            memory_read = 0;
            memory_write = 0;
            branch = 1;
            aluop = 2'b01;
        end
    endcase

end
    
endmodule