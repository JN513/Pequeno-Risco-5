module top (
    input clk
);
    

always @(posedge clk ) begin
    
end

endmodule
